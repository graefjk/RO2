----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.01.2021
-- Design Name: 
-- Module Name: sim_StackU_1_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.env.finish;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sim_StackU_1_tb is
--  Port ( );
end sim_StackU_1_tb;

architecture Behavioral of sim_StackU_1_tb is
component stack
    port(   sPC_i : in std_ulogic_vector(11 downto 0);
            write_or_read_i: in std_ulogic; -- 0 for write, 1 for read
            enable_i: in std_ulogic;
            reset_i: in std_ulogic;
            clk_i: in std_ulogic;
            
            full_o: out std_ulogic;
            empty_o: out std_ulogic;
            
            sStack_o: out std_ulogic_vector(11 downto 0)); 
end component;

signal pc_s: std_ulogic_vector(11 downto 0);
signal write_or_read_s: std_logic;
signal enable_s: std_logic;
signal reset_s: std_logic;
signal clk_s: std_logic;

signal full_s: std_logic;
signal empty_s: std_logic;
signal sStack_s: std_ulogic_vector(11 downto 0);

constant clk_period: time := 20 ns;
constant waitTime: time := 10 ns;

begin

uut: stack port map (
			sPC_i => pc_s, 
			write_or_read_i => write_or_read_s, 
			enable_i => enable_s, 
			reset_i => reset_s, 
			clk_i => clk_s, 
			full_o => full_s, 
			empty_o => empty_s,
			sStack_o => sStack_s);

    clk_process: process
    begin
        clk_s <= '0';
        wait for clk_period / 2;
        clk_s <= '1';
        wait for clk_period / 2;
    end process;
    
	write_or_read_process: process
    begin
        write_or_read_s <= '0';
        wait for 3ns;
        write_or_read_s <= '1';
        wait for 3ns;
    end process;

    
    stimuli: process
    begin
	reset_s <= '0';
	enable_s <= '1';

 wait for waitTime;   
report "The Test has started ";

report "Variant of Stack_tb_long5 with unstable write_or_read_s. ";

wait for waitTime;
pc_s <= "000000000000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000000111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000001111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000010111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000011111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000100111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000101111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000110111";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111000";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111001";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111010";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111011";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111100";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111101";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111110";
wait for waitTime;
wait for waitTime;
pc_s <= "000000111111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001000111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001001111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001010111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001011111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001100111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001101111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110110";
wait for waitTime;
wait for waitTime;
pc_s <= "000001110111";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111000";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111001";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111010";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111011";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111100";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111101";
wait for waitTime;
wait for waitTime;
pc_s <= "000001111110";
wait for waitTime;
wait for waitTime;
pc_s <= "001111001111";
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
wait for waitTime;
report "You can see that this unstable write_or_read_s leads to inconsistency of the Stack ";

report "The Test is finished ";

		finish;
    end process;

end Behavioral;
