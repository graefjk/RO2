		finish;
    end process;

end Behavioral;
