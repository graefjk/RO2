--insert_start_here
--insert_code_here
--insert_end_here
