
    end process;

end Behavioral;
