----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Jannik Graef
-- 
-- Create Date: 04.12.2021 12:00:50
-- Design Name: 
-- Module Name: sim_ALU_tb_LOAD - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sim_ALU_tb_LOAD is
--  Port ( );
end sim_ALU_tb_LOAD;

architecture Behavioral of sim_ALU_tb_LOAD is
component ALU
 Port (sA_i: in std_ulogic_vector(7 downto 0); --input signals
       sB_i: in std_ulogic_vector(7 downto 0);
       opcode_select_i: in std_ulogic_vector(5 downto 0);
       reset_i: in std_logic;
       clk_i: in std_logic;
       enable_i: in std_logic;
       
       sALU_o: out std_ulogic_vector(7 downto 0); -- output signals
       sCARRY_o: out std_logic;
       sZERO_o: out std_logic);
end component;

signal sA_s: std_ulogic_vector(7 downto 0);
signal sB_s: std_ulogic_vector(7 downto 0);
signal opcode_select_s: std_ulogic_vector(5 downto 0);
signal reset_s: std_logic;
signal clk_s: std_logic;
signal enable_s: std_logic;

signal sALU_s: std_ulogic_vector(7 downto 0);
signal sCARRY_s: std_logic;
signal sZERO_s: std_logic;

constant clk_period: time := 20 ns;
constant waitTime: time := 20 ns;

begin

uut: ALU port map (
			sA_i => sA_s,
			sB_i => sB_s,
			opcode_select_i => opcode_select_s, 
			reset_i => reset_s, 
			clk_i => clk_s, 
			enable_i => enable_s,
			sALU_o => sALU_s, 
			sCARRY_o => sCARRY_s, 
			sZERO_o =>sZERO_s);

    clk_process: process
    begin
        clk_s <= '0';
        wait for clk_period / 2;
        clk_s <= '1';
        wait for clk_period / 2;
    end process;
    

    
    stimuli: process
	variable err_cnt: integer := 0; 
    begin
 enable_s <= '1';
 wait for waitTime;   

opcode_select_s <= "001111";sB_s <= "00000000";
wait for waitTime;
assert sALU_s = "00000000"
	report "LOAD error at LOAD 00000000" severity error;

wait for waitTime;
sB_s <= "00000001";
wait for waitTime;
assert sALU_s = "00000001"
	report "LOAD error at LOAD 00000001" severity error;

wait for waitTime;
sB_s <= "00000010";
wait for waitTime;
assert sALU_s = "00000010"
	report "LOAD error at LOAD 00000010" severity error;

wait for waitTime;
sB_s <= "00000011";
wait for waitTime;
assert sALU_s = "00000011"
	report "LOAD error at LOAD 00000011" severity error;

wait for waitTime;
sB_s <= "00000100";
wait for waitTime;
assert sALU_s = "00000100"
	report "LOAD error at LOAD 00000100" severity error;

wait for waitTime;
sB_s <= "00000101";
wait for waitTime;
assert sALU_s = "00000101"
	report "LOAD error at LOAD 00000101" severity error;

wait for waitTime;
sB_s <= "00000110";
wait for waitTime;
assert sALU_s = "00000110"
	report "LOAD error at LOAD 00000110" severity error;

wait for waitTime;
sB_s <= "00000111";
wait for waitTime;
assert sALU_s = "00000111"
	report "LOAD error at LOAD 00000111" severity error;

wait for waitTime;
sB_s <= "00001000";
wait for waitTime;
assert sALU_s = "00001000"
	report "LOAD error at LOAD 00001000" severity error;

wait for waitTime;
sB_s <= "00001001";
wait for waitTime;
assert sALU_s = "00001001"
	report "LOAD error at LOAD 00001001" severity error;

wait for waitTime;
sB_s <= "00001010";
wait for waitTime;
assert sALU_s = "00001010"
	report "LOAD error at LOAD 00001010" severity error;

wait for waitTime;
sB_s <= "00001011";
wait for waitTime;
assert sALU_s = "00001011"
	report "LOAD error at LOAD 00001011" severity error;

wait for waitTime;
sB_s <= "00001100";
wait for waitTime;
assert sALU_s = "00001100"
	report "LOAD error at LOAD 00001100" severity error;

wait for waitTime;
sB_s <= "00001101";
wait for waitTime;
assert sALU_s = "00001101"
	report "LOAD error at LOAD 00001101" severity error;

wait for waitTime;
sB_s <= "00001110";
wait for waitTime;
assert sALU_s = "00001110"
	report "LOAD error at LOAD 00001110" severity error;

wait for waitTime;
sB_s <= "00001111";
wait for waitTime;
assert sALU_s = "00001111"
	report "LOAD error at LOAD 00001111" severity error;

wait for waitTime;
sB_s <= "00010000";
wait for waitTime;
assert sALU_s = "00010000"
	report "LOAD error at LOAD 00010000" severity error;

wait for waitTime;
sB_s <= "00010001";
wait for waitTime;
assert sALU_s = "00010001"
	report "LOAD error at LOAD 00010001" severity error;

wait for waitTime;
sB_s <= "00010010";
wait for waitTime;
assert sALU_s = "00010010"
	report "LOAD error at LOAD 00010010" severity error;

wait for waitTime;
sB_s <= "00010011";
wait for waitTime;
assert sALU_s = "00010011"
	report "LOAD error at LOAD 00010011" severity error;

wait for waitTime;
sB_s <= "00010100";
wait for waitTime;
assert sALU_s = "00010100"
	report "LOAD error at LOAD 00010100" severity error;

wait for waitTime;
sB_s <= "00010101";
wait for waitTime;
assert sALU_s = "00010101"
	report "LOAD error at LOAD 00010101" severity error;

wait for waitTime;
sB_s <= "00010110";
wait for waitTime;
assert sALU_s = "00010110"
	report "LOAD error at LOAD 00010110" severity error;

wait for waitTime;
sB_s <= "00010111";
wait for waitTime;
assert sALU_s = "00010111"
	report "LOAD error at LOAD 00010111" severity error;

wait for waitTime;
sB_s <= "00011000";
wait for waitTime;
assert sALU_s = "00011000"
	report "LOAD error at LOAD 00011000" severity error;

wait for waitTime;
sB_s <= "00011001";
wait for waitTime;
assert sALU_s = "00011001"
	report "LOAD error at LOAD 00011001" severity error;

wait for waitTime;
sB_s <= "00011010";
wait for waitTime;
assert sALU_s = "00011010"
	report "LOAD error at LOAD 00011010" severity error;

wait for waitTime;
sB_s <= "00011011";
wait for waitTime;
assert sALU_s = "00011011"
	report "LOAD error at LOAD 00011011" severity error;

wait for waitTime;
sB_s <= "00011100";
wait for waitTime;
assert sALU_s = "00011100"
	report "LOAD error at LOAD 00011100" severity error;

wait for waitTime;
sB_s <= "00011101";
wait for waitTime;
assert sALU_s = "00011101"
	report "LOAD error at LOAD 00011101" severity error;

wait for waitTime;
sB_s <= "00011110";
wait for waitTime;
assert sALU_s = "00011110"
	report "LOAD error at LOAD 00011110" severity error;

wait for waitTime;
sB_s <= "00011111";
wait for waitTime;
assert sALU_s = "00011111"
	report "LOAD error at LOAD 00011111" severity error;

wait for waitTime;
sB_s <= "00100000";
wait for waitTime;
assert sALU_s = "00100000"
	report "LOAD error at LOAD 00100000" severity error;

wait for waitTime;
sB_s <= "00100001";
wait for waitTime;
assert sALU_s = "00100001"
	report "LOAD error at LOAD 00100001" severity error;

wait for waitTime;
sB_s <= "00100010";
wait for waitTime;
assert sALU_s = "00100010"
	report "LOAD error at LOAD 00100010" severity error;

wait for waitTime;
sB_s <= "00100011";
wait for waitTime;
assert sALU_s = "00100011"
	report "LOAD error at LOAD 00100011" severity error;

wait for waitTime;
sB_s <= "00100100";
wait for waitTime;
assert sALU_s = "00100100"
	report "LOAD error at LOAD 00100100" severity error;

wait for waitTime;
sB_s <= "00100101";
wait for waitTime;
assert sALU_s = "00100101"
	report "LOAD error at LOAD 00100101" severity error;

wait for waitTime;
sB_s <= "00100110";
wait for waitTime;
assert sALU_s = "00100110"
	report "LOAD error at LOAD 00100110" severity error;

wait for waitTime;
sB_s <= "00100111";
wait for waitTime;
assert sALU_s = "00100111"
	report "LOAD error at LOAD 00100111" severity error;

wait for waitTime;
sB_s <= "00101000";
wait for waitTime;
assert sALU_s = "00101000"
	report "LOAD error at LOAD 00101000" severity error;

wait for waitTime;
sB_s <= "00101001";
wait for waitTime;
assert sALU_s = "00101001"
	report "LOAD error at LOAD 00101001" severity error;

wait for waitTime;
sB_s <= "00101010";
wait for waitTime;
assert sALU_s = "00101010"
	report "LOAD error at LOAD 00101010" severity error;

wait for waitTime;
sB_s <= "00101011";
wait for waitTime;
assert sALU_s = "00101011"
	report "LOAD error at LOAD 00101011" severity error;

wait for waitTime;
sB_s <= "00101100";
wait for waitTime;
assert sALU_s = "00101100"
	report "LOAD error at LOAD 00101100" severity error;

wait for waitTime;
sB_s <= "00101101";
wait for waitTime;
assert sALU_s = "00101101"
	report "LOAD error at LOAD 00101101" severity error;

wait for waitTime;
sB_s <= "00101110";
wait for waitTime;
assert sALU_s = "00101110"
	report "LOAD error at LOAD 00101110" severity error;

wait for waitTime;
sB_s <= "00101111";
wait for waitTime;
assert sALU_s = "00101111"
	report "LOAD error at LOAD 00101111" severity error;

wait for waitTime;
sB_s <= "00110000";
wait for waitTime;
assert sALU_s = "00110000"
	report "LOAD error at LOAD 00110000" severity error;

wait for waitTime;
sB_s <= "00110001";
wait for waitTime;
assert sALU_s = "00110001"
	report "LOAD error at LOAD 00110001" severity error;

wait for waitTime;
sB_s <= "00110010";
wait for waitTime;
assert sALU_s = "00110010"
	report "LOAD error at LOAD 00110010" severity error;

wait for waitTime;
sB_s <= "00110011";
wait for waitTime;
assert sALU_s = "00110011"
	report "LOAD error at LOAD 00110011" severity error;

wait for waitTime;
sB_s <= "00110100";
wait for waitTime;
assert sALU_s = "00110100"
	report "LOAD error at LOAD 00110100" severity error;

wait for waitTime;
sB_s <= "00110101";
wait for waitTime;
assert sALU_s = "00110101"
	report "LOAD error at LOAD 00110101" severity error;

wait for waitTime;
sB_s <= "00110110";
wait for waitTime;
assert sALU_s = "00110110"
	report "LOAD error at LOAD 00110110" severity error;

wait for waitTime;
sB_s <= "00110111";
wait for waitTime;
assert sALU_s = "00110111"
	report "LOAD error at LOAD 00110111" severity error;

wait for waitTime;
sB_s <= "00111000";
wait for waitTime;
assert sALU_s = "00111000"
	report "LOAD error at LOAD 00111000" severity error;

wait for waitTime;
sB_s <= "00111001";
wait for waitTime;
assert sALU_s = "00111001"
	report "LOAD error at LOAD 00111001" severity error;

wait for waitTime;
sB_s <= "00111010";
wait for waitTime;
assert sALU_s = "00111010"
	report "LOAD error at LOAD 00111010" severity error;

wait for waitTime;
sB_s <= "00111011";
wait for waitTime;
assert sALU_s = "00111011"
	report "LOAD error at LOAD 00111011" severity error;

wait for waitTime;
sB_s <= "00111100";
wait for waitTime;
assert sALU_s = "00111100"
	report "LOAD error at LOAD 00111100" severity error;

wait for waitTime;
sB_s <= "00111101";
wait for waitTime;
assert sALU_s = "00111101"
	report "LOAD error at LOAD 00111101" severity error;

wait for waitTime;
sB_s <= "00111110";
wait for waitTime;
assert sALU_s = "00111110"
	report "LOAD error at LOAD 00111110" severity error;

wait for waitTime;
sB_s <= "00111111";
wait for waitTime;
assert sALU_s = "00111111"
	report "LOAD error at LOAD 00111111" severity error;

wait for waitTime;
sB_s <= "01000000";
wait for waitTime;
assert sALU_s = "01000000"
	report "LOAD error at LOAD 01000000" severity error;

wait for waitTime;
sB_s <= "01000001";
wait for waitTime;
assert sALU_s = "01000001"
	report "LOAD error at LOAD 01000001" severity error;

wait for waitTime;
sB_s <= "01000010";
wait for waitTime;
assert sALU_s = "01000010"
	report "LOAD error at LOAD 01000010" severity error;

wait for waitTime;
sB_s <= "01000011";
wait for waitTime;
assert sALU_s = "01000011"
	report "LOAD error at LOAD 01000011" severity error;

wait for waitTime;
sB_s <= "01000100";
wait for waitTime;
assert sALU_s = "01000100"
	report "LOAD error at LOAD 01000100" severity error;

wait for waitTime;
sB_s <= "01000101";
wait for waitTime;
assert sALU_s = "01000101"
	report "LOAD error at LOAD 01000101" severity error;

wait for waitTime;
sB_s <= "01000110";
wait for waitTime;
assert sALU_s = "01000110"
	report "LOAD error at LOAD 01000110" severity error;

wait for waitTime;
sB_s <= "01000111";
wait for waitTime;
assert sALU_s = "01000111"
	report "LOAD error at LOAD 01000111" severity error;

wait for waitTime;
sB_s <= "01001000";
wait for waitTime;
assert sALU_s = "01001000"
	report "LOAD error at LOAD 01001000" severity error;

wait for waitTime;
sB_s <= "01001001";
wait for waitTime;
assert sALU_s = "01001001"
	report "LOAD error at LOAD 01001001" severity error;

wait for waitTime;
sB_s <= "01001010";
wait for waitTime;
assert sALU_s = "01001010"
	report "LOAD error at LOAD 01001010" severity error;

wait for waitTime;
sB_s <= "01001011";
wait for waitTime;
assert sALU_s = "01001011"
	report "LOAD error at LOAD 01001011" severity error;

wait for waitTime;
sB_s <= "01001100";
wait for waitTime;
assert sALU_s = "01001100"
	report "LOAD error at LOAD 01001100" severity error;

wait for waitTime;
sB_s <= "01001101";
wait for waitTime;
assert sALU_s = "01001101"
	report "LOAD error at LOAD 01001101" severity error;

wait for waitTime;
sB_s <= "01001110";
wait for waitTime;
assert sALU_s = "01001110"
	report "LOAD error at LOAD 01001110" severity error;

wait for waitTime;
sB_s <= "01001111";
wait for waitTime;
assert sALU_s = "01001111"
	report "LOAD error at LOAD 01001111" severity error;

wait for waitTime;
sB_s <= "01010000";
wait for waitTime;
assert sALU_s = "01010000"
	report "LOAD error at LOAD 01010000" severity error;

wait for waitTime;
sB_s <= "01010001";
wait for waitTime;
assert sALU_s = "01010001"
	report "LOAD error at LOAD 01010001" severity error;

wait for waitTime;
sB_s <= "01010010";
wait for waitTime;
assert sALU_s = "01010010"
	report "LOAD error at LOAD 01010010" severity error;

wait for waitTime;
sB_s <= "01010011";
wait for waitTime;
assert sALU_s = "01010011"
	report "LOAD error at LOAD 01010011" severity error;

wait for waitTime;
sB_s <= "01010100";
wait for waitTime;
assert sALU_s = "01010100"
	report "LOAD error at LOAD 01010100" severity error;

wait for waitTime;
sB_s <= "01010101";
wait for waitTime;
assert sALU_s = "01010101"
	report "LOAD error at LOAD 01010101" severity error;

wait for waitTime;
sB_s <= "01010110";
wait for waitTime;
assert sALU_s = "01010110"
	report "LOAD error at LOAD 01010110" severity error;

wait for waitTime;
sB_s <= "01010111";
wait for waitTime;
assert sALU_s = "01010111"
	report "LOAD error at LOAD 01010111" severity error;

wait for waitTime;
sB_s <= "01011000";
wait for waitTime;
assert sALU_s = "01011000"
	report "LOAD error at LOAD 01011000" severity error;

wait for waitTime;
sB_s <= "01011001";
wait for waitTime;
assert sALU_s = "01011001"
	report "LOAD error at LOAD 01011001" severity error;

wait for waitTime;
sB_s <= "01011010";
wait for waitTime;
assert sALU_s = "01011010"
	report "LOAD error at LOAD 01011010" severity error;

wait for waitTime;
sB_s <= "01011011";
wait for waitTime;
assert sALU_s = "01011011"
	report "LOAD error at LOAD 01011011" severity error;

wait for waitTime;
sB_s <= "01011100";
wait for waitTime;
assert sALU_s = "01011100"
	report "LOAD error at LOAD 01011100" severity error;

wait for waitTime;
sB_s <= "01011101";
wait for waitTime;
assert sALU_s = "01011101"
	report "LOAD error at LOAD 01011101" severity error;

wait for waitTime;
sB_s <= "01011110";
wait for waitTime;
assert sALU_s = "01011110"
	report "LOAD error at LOAD 01011110" severity error;

wait for waitTime;
sB_s <= "01011111";
wait for waitTime;
assert sALU_s = "01011111"
	report "LOAD error at LOAD 01011111" severity error;

wait for waitTime;
sB_s <= "01100000";
wait for waitTime;
assert sALU_s = "01100000"
	report "LOAD error at LOAD 01100000" severity error;

wait for waitTime;
sB_s <= "01100001";
wait for waitTime;
assert sALU_s = "01100001"
	report "LOAD error at LOAD 01100001" severity error;

wait for waitTime;
sB_s <= "01100010";
wait for waitTime;
assert sALU_s = "01100010"
	report "LOAD error at LOAD 01100010" severity error;

wait for waitTime;
sB_s <= "01100011";
wait for waitTime;
assert sALU_s = "01100011"
	report "LOAD error at LOAD 01100011" severity error;

wait for waitTime;
sB_s <= "01100100";
wait for waitTime;
assert sALU_s = "01100100"
	report "LOAD error at LOAD 01100100" severity error;

wait for waitTime;
sB_s <= "01100101";
wait for waitTime;
assert sALU_s = "01100101"
	report "LOAD error at LOAD 01100101" severity error;

wait for waitTime;
sB_s <= "01100110";
wait for waitTime;
assert sALU_s = "01100110"
	report "LOAD error at LOAD 01100110" severity error;

wait for waitTime;
sB_s <= "01100111";
wait for waitTime;
assert sALU_s = "01100111"
	report "LOAD error at LOAD 01100111" severity error;

wait for waitTime;
sB_s <= "01101000";
wait for waitTime;
assert sALU_s = "01101000"
	report "LOAD error at LOAD 01101000" severity error;

wait for waitTime;
sB_s <= "01101001";
wait for waitTime;
assert sALU_s = "01101001"
	report "LOAD error at LOAD 01101001" severity error;

wait for waitTime;
sB_s <= "01101010";
wait for waitTime;
assert sALU_s = "01101010"
	report "LOAD error at LOAD 01101010" severity error;

wait for waitTime;
sB_s <= "01101011";
wait for waitTime;
assert sALU_s = "01101011"
	report "LOAD error at LOAD 01101011" severity error;

wait for waitTime;
sB_s <= "01101100";
wait for waitTime;
assert sALU_s = "01101100"
	report "LOAD error at LOAD 01101100" severity error;

wait for waitTime;
sB_s <= "01101101";
wait for waitTime;
assert sALU_s = "01101101"
	report "LOAD error at LOAD 01101101" severity error;

wait for waitTime;
sB_s <= "01101110";
wait for waitTime;
assert sALU_s = "01101110"
	report "LOAD error at LOAD 01101110" severity error;

wait for waitTime;
sB_s <= "01101111";
wait for waitTime;
assert sALU_s = "01101111"
	report "LOAD error at LOAD 01101111" severity error;

wait for waitTime;
sB_s <= "01110000";
wait for waitTime;
assert sALU_s = "01110000"
	report "LOAD error at LOAD 01110000" severity error;

wait for waitTime;
sB_s <= "01110001";
wait for waitTime;
assert sALU_s = "01110001"
	report "LOAD error at LOAD 01110001" severity error;

wait for waitTime;
sB_s <= "01110010";
wait for waitTime;
assert sALU_s = "01110010"
	report "LOAD error at LOAD 01110010" severity error;

wait for waitTime;
sB_s <= "01110011";
wait for waitTime;
assert sALU_s = "01110011"
	report "LOAD error at LOAD 01110011" severity error;

wait for waitTime;
sB_s <= "01110100";
wait for waitTime;
assert sALU_s = "01110100"
	report "LOAD error at LOAD 01110100" severity error;

wait for waitTime;
sB_s <= "01110101";
wait for waitTime;
assert sALU_s = "01110101"
	report "LOAD error at LOAD 01110101" severity error;

wait for waitTime;
sB_s <= "01110110";
wait for waitTime;
assert sALU_s = "01110110"
	report "LOAD error at LOAD 01110110" severity error;

wait for waitTime;
sB_s <= "01110111";
wait for waitTime;
assert sALU_s = "01110111"
	report "LOAD error at LOAD 01110111" severity error;

wait for waitTime;
sB_s <= "01111000";
wait for waitTime;
assert sALU_s = "01111000"
	report "LOAD error at LOAD 01111000" severity error;

wait for waitTime;
sB_s <= "01111001";
wait for waitTime;
assert sALU_s = "01111001"
	report "LOAD error at LOAD 01111001" severity error;

wait for waitTime;
sB_s <= "01111010";
wait for waitTime;
assert sALU_s = "01111010"
	report "LOAD error at LOAD 01111010" severity error;

wait for waitTime;
sB_s <= "01111011";
wait for waitTime;
assert sALU_s = "01111011"
	report "LOAD error at LOAD 01111011" severity error;

wait for waitTime;
sB_s <= "01111100";
wait for waitTime;
assert sALU_s = "01111100"
	report "LOAD error at LOAD 01111100" severity error;

wait for waitTime;
sB_s <= "01111101";
wait for waitTime;
assert sALU_s = "01111101"
	report "LOAD error at LOAD 01111101" severity error;

wait for waitTime;
sB_s <= "01111110";
wait for waitTime;
assert sALU_s = "01111110"
	report "LOAD error at LOAD 01111110" severity error;

wait for waitTime;
sB_s <= "01111111";
wait for waitTime;
assert sALU_s = "01111111"
	report "LOAD error at LOAD 01111111" severity error;

wait for waitTime;
sB_s <= "10000000";
wait for waitTime;
assert sALU_s = "10000000"
	report "LOAD error at LOAD 10000000" severity error;

wait for waitTime;
sB_s <= "10000001";
wait for waitTime;
assert sALU_s = "10000001"
	report "LOAD error at LOAD 10000001" severity error;

wait for waitTime;
sB_s <= "10000010";
wait for waitTime;
assert sALU_s = "10000010"
	report "LOAD error at LOAD 10000010" severity error;

wait for waitTime;
sB_s <= "10000011";
wait for waitTime;
assert sALU_s = "10000011"
	report "LOAD error at LOAD 10000011" severity error;

wait for waitTime;
sB_s <= "10000100";
wait for waitTime;
assert sALU_s = "10000100"
	report "LOAD error at LOAD 10000100" severity error;

wait for waitTime;
sB_s <= "10000101";
wait for waitTime;
assert sALU_s = "10000101"
	report "LOAD error at LOAD 10000101" severity error;

wait for waitTime;
sB_s <= "10000110";
wait for waitTime;
assert sALU_s = "10000110"
	report "LOAD error at LOAD 10000110" severity error;

wait for waitTime;
sB_s <= "10000111";
wait for waitTime;
assert sALU_s = "10000111"
	report "LOAD error at LOAD 10000111" severity error;

wait for waitTime;
sB_s <= "10001000";
wait for waitTime;
assert sALU_s = "10001000"
	report "LOAD error at LOAD 10001000" severity error;

wait for waitTime;
sB_s <= "10001001";
wait for waitTime;
assert sALU_s = "10001001"
	report "LOAD error at LOAD 10001001" severity error;

wait for waitTime;
sB_s <= "10001010";
wait for waitTime;
assert sALU_s = "10001010"
	report "LOAD error at LOAD 10001010" severity error;

wait for waitTime;
sB_s <= "10001011";
wait for waitTime;
assert sALU_s = "10001011"
	report "LOAD error at LOAD 10001011" severity error;

wait for waitTime;
sB_s <= "10001100";
wait for waitTime;
assert sALU_s = "10001100"
	report "LOAD error at LOAD 10001100" severity error;

wait for waitTime;
sB_s <= "10001101";
wait for waitTime;
assert sALU_s = "10001101"
	report "LOAD error at LOAD 10001101" severity error;

wait for waitTime;
sB_s <= "10001110";
wait for waitTime;
assert sALU_s = "10001110"
	report "LOAD error at LOAD 10001110" severity error;

wait for waitTime;
sB_s <= "10001111";
wait for waitTime;
assert sALU_s = "10001111"
	report "LOAD error at LOAD 10001111" severity error;

wait for waitTime;
sB_s <= "10010000";
wait for waitTime;
assert sALU_s = "10010000"
	report "LOAD error at LOAD 10010000" severity error;

wait for waitTime;
sB_s <= "10010001";
wait for waitTime;
assert sALU_s = "10010001"
	report "LOAD error at LOAD 10010001" severity error;

wait for waitTime;
sB_s <= "10010010";
wait for waitTime;
assert sALU_s = "10010010"
	report "LOAD error at LOAD 10010010" severity error;

wait for waitTime;
sB_s <= "10010011";
wait for waitTime;
assert sALU_s = "10010011"
	report "LOAD error at LOAD 10010011" severity error;

wait for waitTime;
sB_s <= "10010100";
wait for waitTime;
assert sALU_s = "10010100"
	report "LOAD error at LOAD 10010100" severity error;

wait for waitTime;
sB_s <= "10010101";
wait for waitTime;
assert sALU_s = "10010101"
	report "LOAD error at LOAD 10010101" severity error;

wait for waitTime;
sB_s <= "10010110";
wait for waitTime;
assert sALU_s = "10010110"
	report "LOAD error at LOAD 10010110" severity error;

wait for waitTime;
sB_s <= "10010111";
wait for waitTime;
assert sALU_s = "10010111"
	report "LOAD error at LOAD 10010111" severity error;

wait for waitTime;
sB_s <= "10011000";
wait for waitTime;
assert sALU_s = "10011000"
	report "LOAD error at LOAD 10011000" severity error;

wait for waitTime;
sB_s <= "10011001";
wait for waitTime;
assert sALU_s = "10011001"
	report "LOAD error at LOAD 10011001" severity error;

wait for waitTime;
sB_s <= "10011010";
wait for waitTime;
assert sALU_s = "10011010"
	report "LOAD error at LOAD 10011010" severity error;

wait for waitTime;
sB_s <= "10011011";
wait for waitTime;
assert sALU_s = "10011011"
	report "LOAD error at LOAD 10011011" severity error;

wait for waitTime;
sB_s <= "10011100";
wait for waitTime;
assert sALU_s = "10011100"
	report "LOAD error at LOAD 10011100" severity error;

wait for waitTime;
sB_s <= "10011101";
wait for waitTime;
assert sALU_s = "10011101"
	report "LOAD error at LOAD 10011101" severity error;

wait for waitTime;
sB_s <= "10011110";
wait for waitTime;
assert sALU_s = "10011110"
	report "LOAD error at LOAD 10011110" severity error;

wait for waitTime;
sB_s <= "10011111";
wait for waitTime;
assert sALU_s = "10011111"
	report "LOAD error at LOAD 10011111" severity error;

wait for waitTime;
sB_s <= "10100000";
wait for waitTime;
assert sALU_s = "10100000"
	report "LOAD error at LOAD 10100000" severity error;

wait for waitTime;
sB_s <= "10100001";
wait for waitTime;
assert sALU_s = "10100001"
	report "LOAD error at LOAD 10100001" severity error;

wait for waitTime;
sB_s <= "10100010";
wait for waitTime;
assert sALU_s = "10100010"
	report "LOAD error at LOAD 10100010" severity error;

wait for waitTime;
sB_s <= "10100011";
wait for waitTime;
assert sALU_s = "10100011"
	report "LOAD error at LOAD 10100011" severity error;

wait for waitTime;
sB_s <= "10100100";
wait for waitTime;
assert sALU_s = "10100100"
	report "LOAD error at LOAD 10100100" severity error;

wait for waitTime;
sB_s <= "10100101";
wait for waitTime;
assert sALU_s = "10100101"
	report "LOAD error at LOAD 10100101" severity error;

wait for waitTime;
sB_s <= "10100110";
wait for waitTime;
assert sALU_s = "10100110"
	report "LOAD error at LOAD 10100110" severity error;

wait for waitTime;
sB_s <= "10100111";
wait for waitTime;
assert sALU_s = "10100111"
	report "LOAD error at LOAD 10100111" severity error;

wait for waitTime;
sB_s <= "10101000";
wait for waitTime;
assert sALU_s = "10101000"
	report "LOAD error at LOAD 10101000" severity error;

wait for waitTime;
sB_s <= "10101001";
wait for waitTime;
assert sALU_s = "10101001"
	report "LOAD error at LOAD 10101001" severity error;

wait for waitTime;
sB_s <= "10101010";
wait for waitTime;
assert sALU_s = "10101010"
	report "LOAD error at LOAD 10101010" severity error;

wait for waitTime;
sB_s <= "10101011";
wait for waitTime;
assert sALU_s = "10101011"
	report "LOAD error at LOAD 10101011" severity error;

wait for waitTime;
sB_s <= "10101100";
wait for waitTime;
assert sALU_s = "10101100"
	report "LOAD error at LOAD 10101100" severity error;

wait for waitTime;
sB_s <= "10101101";
wait for waitTime;
assert sALU_s = "10101101"
	report "LOAD error at LOAD 10101101" severity error;

wait for waitTime;
sB_s <= "10101110";
wait for waitTime;
assert sALU_s = "10101110"
	report "LOAD error at LOAD 10101110" severity error;

wait for waitTime;
sB_s <= "10101111";
wait for waitTime;
assert sALU_s = "10101111"
	report "LOAD error at LOAD 10101111" severity error;

wait for waitTime;
sB_s <= "10110000";
wait for waitTime;
assert sALU_s = "10110000"
	report "LOAD error at LOAD 10110000" severity error;

wait for waitTime;
sB_s <= "10110001";
wait for waitTime;
assert sALU_s = "10110001"
	report "LOAD error at LOAD 10110001" severity error;

wait for waitTime;
sB_s <= "10110010";
wait for waitTime;
assert sALU_s = "10110010"
	report "LOAD error at LOAD 10110010" severity error;

wait for waitTime;
sB_s <= "10110011";
wait for waitTime;
assert sALU_s = "10110011"
	report "LOAD error at LOAD 10110011" severity error;

wait for waitTime;
sB_s <= "10110100";
wait for waitTime;
assert sALU_s = "10110100"
	report "LOAD error at LOAD 10110100" severity error;

wait for waitTime;
sB_s <= "10110101";
wait for waitTime;
assert sALU_s = "10110101"
	report "LOAD error at LOAD 10110101" severity error;

wait for waitTime;
sB_s <= "10110110";
wait for waitTime;
assert sALU_s = "10110110"
	report "LOAD error at LOAD 10110110" severity error;

wait for waitTime;
sB_s <= "10110111";
wait for waitTime;
assert sALU_s = "10110111"
	report "LOAD error at LOAD 10110111" severity error;

wait for waitTime;
sB_s <= "10111000";
wait for waitTime;
assert sALU_s = "10111000"
	report "LOAD error at LOAD 10111000" severity error;

wait for waitTime;
sB_s <= "10111001";
wait for waitTime;
assert sALU_s = "10111001"
	report "LOAD error at LOAD 10111001" severity error;

wait for waitTime;
sB_s <= "10111010";
wait for waitTime;
assert sALU_s = "10111010"
	report "LOAD error at LOAD 10111010" severity error;

wait for waitTime;
sB_s <= "10111011";
wait for waitTime;
assert sALU_s = "10111011"
	report "LOAD error at LOAD 10111011" severity error;

wait for waitTime;
sB_s <= "10111100";
wait for waitTime;
assert sALU_s = "10111100"
	report "LOAD error at LOAD 10111100" severity error;

wait for waitTime;
sB_s <= "10111101";
wait for waitTime;
assert sALU_s = "10111101"
	report "LOAD error at LOAD 10111101" severity error;

wait for waitTime;
sB_s <= "10111110";
wait for waitTime;
assert sALU_s = "10111110"
	report "LOAD error at LOAD 10111110" severity error;

wait for waitTime;
sB_s <= "10111111";
wait for waitTime;
assert sALU_s = "10111111"
	report "LOAD error at LOAD 10111111" severity error;

wait for waitTime;
sB_s <= "11000000";
wait for waitTime;
assert sALU_s = "11000000"
	report "LOAD error at LOAD 11000000" severity error;

wait for waitTime;
sB_s <= "11000001";
wait for waitTime;
assert sALU_s = "11000001"
	report "LOAD error at LOAD 11000001" severity error;

wait for waitTime;
sB_s <= "11000010";
wait for waitTime;
assert sALU_s = "11000010"
	report "LOAD error at LOAD 11000010" severity error;

wait for waitTime;
sB_s <= "11000011";
wait for waitTime;
assert sALU_s = "11000011"
	report "LOAD error at LOAD 11000011" severity error;

wait for waitTime;
sB_s <= "11000100";
wait for waitTime;
assert sALU_s = "11000100"
	report "LOAD error at LOAD 11000100" severity error;

wait for waitTime;
sB_s <= "11000101";
wait for waitTime;
assert sALU_s = "11000101"
	report "LOAD error at LOAD 11000101" severity error;

wait for waitTime;
sB_s <= "11000110";
wait for waitTime;
assert sALU_s = "11000110"
	report "LOAD error at LOAD 11000110" severity error;

wait for waitTime;
sB_s <= "11000111";
wait for waitTime;
assert sALU_s = "11000111"
	report "LOAD error at LOAD 11000111" severity error;

wait for waitTime;
sB_s <= "11001000";
wait for waitTime;
assert sALU_s = "11001000"
	report "LOAD error at LOAD 11001000" severity error;

wait for waitTime;
sB_s <= "11001001";
wait for waitTime;
assert sALU_s = "11001001"
	report "LOAD error at LOAD 11001001" severity error;

wait for waitTime;
sB_s <= "11001010";
wait for waitTime;
assert sALU_s = "11001010"
	report "LOAD error at LOAD 11001010" severity error;

wait for waitTime;
sB_s <= "11001011";
wait for waitTime;
assert sALU_s = "11001011"
	report "LOAD error at LOAD 11001011" severity error;

wait for waitTime;
sB_s <= "11001100";
wait for waitTime;
assert sALU_s = "11001100"
	report "LOAD error at LOAD 11001100" severity error;

wait for waitTime;
sB_s <= "11001101";
wait for waitTime;
assert sALU_s = "11001101"
	report "LOAD error at LOAD 11001101" severity error;

wait for waitTime;
sB_s <= "11001110";
wait for waitTime;
assert sALU_s = "11001110"
	report "LOAD error at LOAD 11001110" severity error;

wait for waitTime;
sB_s <= "11001111";
wait for waitTime;
assert sALU_s = "11001111"
	report "LOAD error at LOAD 11001111" severity error;

wait for waitTime;
sB_s <= "11010000";
wait for waitTime;
assert sALU_s = "11010000"
	report "LOAD error at LOAD 11010000" severity error;

wait for waitTime;
sB_s <= "11010001";
wait for waitTime;
assert sALU_s = "11010001"
	report "LOAD error at LOAD 11010001" severity error;

wait for waitTime;
sB_s <= "11010010";
wait for waitTime;
assert sALU_s = "11010010"
	report "LOAD error at LOAD 11010010" severity error;

wait for waitTime;
sB_s <= "11010011";
wait for waitTime;
assert sALU_s = "11010011"
	report "LOAD error at LOAD 11010011" severity error;

wait for waitTime;
sB_s <= "11010100";
wait for waitTime;
assert sALU_s = "11010100"
	report "LOAD error at LOAD 11010100" severity error;

wait for waitTime;
sB_s <= "11010101";
wait for waitTime;
assert sALU_s = "11010101"
	report "LOAD error at LOAD 11010101" severity error;

wait for waitTime;
sB_s <= "11010110";
wait for waitTime;
assert sALU_s = "11010110"
	report "LOAD error at LOAD 11010110" severity error;

wait for waitTime;
sB_s <= "11010111";
wait for waitTime;
assert sALU_s = "11010111"
	report "LOAD error at LOAD 11010111" severity error;

wait for waitTime;
sB_s <= "11011000";
wait for waitTime;
assert sALU_s = "11011000"
	report "LOAD error at LOAD 11011000" severity error;

wait for waitTime;
sB_s <= "11011001";
wait for waitTime;
assert sALU_s = "11011001"
	report "LOAD error at LOAD 11011001" severity error;

wait for waitTime;
sB_s <= "11011010";
wait for waitTime;
assert sALU_s = "11011010"
	report "LOAD error at LOAD 11011010" severity error;

wait for waitTime;
sB_s <= "11011011";
wait for waitTime;
assert sALU_s = "11011011"
	report "LOAD error at LOAD 11011011" severity error;

wait for waitTime;
sB_s <= "11011100";
wait for waitTime;
assert sALU_s = "11011100"
	report "LOAD error at LOAD 11011100" severity error;

wait for waitTime;
sB_s <= "11011101";
wait for waitTime;
assert sALU_s = "11011101"
	report "LOAD error at LOAD 11011101" severity error;

wait for waitTime;
sB_s <= "11011110";
wait for waitTime;
assert sALU_s = "11011110"
	report "LOAD error at LOAD 11011110" severity error;

wait for waitTime;
sB_s <= "11011111";
wait for waitTime;
assert sALU_s = "11011111"
	report "LOAD error at LOAD 11011111" severity error;

wait for waitTime;
sB_s <= "11100000";
wait for waitTime;
assert sALU_s = "11100000"
	report "LOAD error at LOAD 11100000" severity error;

wait for waitTime;
sB_s <= "11100001";
wait for waitTime;
assert sALU_s = "11100001"
	report "LOAD error at LOAD 11100001" severity error;

wait for waitTime;
sB_s <= "11100010";
wait for waitTime;
assert sALU_s = "11100010"
	report "LOAD error at LOAD 11100010" severity error;

wait for waitTime;
sB_s <= "11100011";
wait for waitTime;
assert sALU_s = "11100011"
	report "LOAD error at LOAD 11100011" severity error;

wait for waitTime;
sB_s <= "11100100";
wait for waitTime;
assert sALU_s = "11100100"
	report "LOAD error at LOAD 11100100" severity error;

wait for waitTime;
sB_s <= "11100101";
wait for waitTime;
assert sALU_s = "11100101"
	report "LOAD error at LOAD 11100101" severity error;

wait for waitTime;
sB_s <= "11100110";
wait for waitTime;
assert sALU_s = "11100110"
	report "LOAD error at LOAD 11100110" severity error;

wait for waitTime;
sB_s <= "11100111";
wait for waitTime;
assert sALU_s = "11100111"
	report "LOAD error at LOAD 11100111" severity error;

wait for waitTime;
sB_s <= "11101000";
wait for waitTime;
assert sALU_s = "11101000"
	report "LOAD error at LOAD 11101000" severity error;

wait for waitTime;
sB_s <= "11101001";
wait for waitTime;
assert sALU_s = "11101001"
	report "LOAD error at LOAD 11101001" severity error;

wait for waitTime;
sB_s <= "11101010";
wait for waitTime;
assert sALU_s = "11101010"
	report "LOAD error at LOAD 11101010" severity error;

wait for waitTime;
sB_s <= "11101011";
wait for waitTime;
assert sALU_s = "11101011"
	report "LOAD error at LOAD 11101011" severity error;

wait for waitTime;
sB_s <= "11101100";
wait for waitTime;
assert sALU_s = "11101100"
	report "LOAD error at LOAD 11101100" severity error;

wait for waitTime;
sB_s <= "11101101";
wait for waitTime;
assert sALU_s = "11101101"
	report "LOAD error at LOAD 11101101" severity error;

wait for waitTime;
sB_s <= "11101110";
wait for waitTime;
assert sALU_s = "11101110"
	report "LOAD error at LOAD 11101110" severity error;

wait for waitTime;
sB_s <= "11101111";
wait for waitTime;
assert sALU_s = "11101111"
	report "LOAD error at LOAD 11101111" severity error;

wait for waitTime;
sB_s <= "11110000";
wait for waitTime;
assert sALU_s = "11110000"
	report "LOAD error at LOAD 11110000" severity error;

wait for waitTime;
sB_s <= "11110001";
wait for waitTime;
assert sALU_s = "11110001"
	report "LOAD error at LOAD 11110001" severity error;

wait for waitTime;
sB_s <= "11110010";
wait for waitTime;
assert sALU_s = "11110010"
	report "LOAD error at LOAD 11110010" severity error;

wait for waitTime;
sB_s <= "11110011";
wait for waitTime;
assert sALU_s = "11110011"
	report "LOAD error at LOAD 11110011" severity error;

wait for waitTime;
sB_s <= "11110100";
wait for waitTime;
assert sALU_s = "11110100"
	report "LOAD error at LOAD 11110100" severity error;

wait for waitTime;
sB_s <= "11110101";
wait for waitTime;
assert sALU_s = "11110101"
	report "LOAD error at LOAD 11110101" severity error;

wait for waitTime;
sB_s <= "11110110";
wait for waitTime;
assert sALU_s = "11110110"
	report "LOAD error at LOAD 11110110" severity error;

wait for waitTime;
sB_s <= "11110111";
wait for waitTime;
assert sALU_s = "11110111"
	report "LOAD error at LOAD 11110111" severity error;

wait for waitTime;
sB_s <= "11111000";
wait for waitTime;
assert sALU_s = "11111000"
	report "LOAD error at LOAD 11111000" severity error;

wait for waitTime;
sB_s <= "11111001";
wait for waitTime;
assert sALU_s = "11111001"
	report "LOAD error at LOAD 11111001" severity error;

wait for waitTime;
sB_s <= "11111010";
wait for waitTime;
assert sALU_s = "11111010"
	report "LOAD error at LOAD 11111010" severity error;

wait for waitTime;
sB_s <= "11111011";
wait for waitTime;
assert sALU_s = "11111011"
	report "LOAD error at LOAD 11111011" severity error;

wait for waitTime;
sB_s <= "11111100";
wait for waitTime;
assert sALU_s = "11111100"
	report "LOAD error at LOAD 11111100" severity error;

wait for waitTime;
sB_s <= "11111101";
wait for waitTime;
assert sALU_s = "11111101"
	report "LOAD error at LOAD 11111101" severity error;

wait for waitTime;
sB_s <= "11111110";
wait for waitTime;
assert sALU_s = "11111110"
	report "LOAD error at LOAD 11111110" severity error;

wait for waitTime;
sB_s <= "11111111";
wait for waitTime;
assert sALU_s = "11111111"
	report "LOAD error at LOAD 11111111" severity error;

wait for waitTime;


    end process;

end Behavioral;
