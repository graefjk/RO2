--insert_code_here
